module tb_render();
	import video_types::*;
	 initial $display("work dammit");

endmodule
