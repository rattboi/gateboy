/*
* Project: Gateboy
*
*
*/

module testbench;


always begin
    $display("Hello Testbench");
    $finish;
end

endmodule
