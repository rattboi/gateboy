/* Project: Gateboy
 * Authors: Tyler Tricker
 * 
 * Description: testbench
 */
 
 module testbench;
 
 always
  begin
     $display("Hello Test Benched World");
	  $finish();
  end
 
 endmodule
 