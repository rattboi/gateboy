module tb_render();
	import video_types::*;
	$display("work dammit");

endmodule
