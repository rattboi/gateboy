module tb_render();


endmodule
